timeunit 1us/100ns;

// this is a comment
module top;
  // this is another comment
  initial begin
    $display("hello, world!");
  end // end module top
endmodule
